//=======================================================================
// COPYRIGHT (C) 2018-2020 RockerIC, Ltd.
// This software and the associated documentation are confidential and
// proprietary to RockerIC, Ltd. Your use or disclosure of this software
// is subject to the terms and conditions of a consulting agreement
// between you, or your company, and RockerIC, Ltd. In the event of
// publications, the following notice is applicable:
//
// ALL RIGHTS RESERVED
//
// The entire notice above must be reproduced on all authorized copies.
//
// VisitUs  : www.rockeric.com
// Support  : support@rockeric.com
// WeChat   : eva_bill
//-----------------------------------------------------------------------
`ifndef LVC_I2C_MONITOR_COMMON_SV
`define LVC_I2C_MONITOR_COMMON_SV

typedef class lvc_i2c_master_transaction;
typedef class lvc_i2c_slave_transaction;

class lvc_i2c_monitor_common extends uvm_object;

  lvc_i2c_vif i2c_if;
  lvc_i2c_agent_configuration cfg;

  logic   trans_start_flag = 0;
  logic   trans_stop_flag = 0;
  logic   trans_restart_flag = 0;
  int unsigned ack_count=0;  //count ack
  int unsigned nack_count=0;  //count nak
  bit[7:0] mon_data[$];
  int mon_data_index = 0;
  `uvm_object_utils_begin(lvc_i2c_monitor_common)
  `uvm_object_utils_end

  function new(string name = "lvc_i2c_monitor_common");
    super.new(name);
  endfunction

  extern virtual function void assign_vif(lvc_i2c_vif i2c_if);
  extern virtual task source_event(event sv_e, uvm_event uvm_e);
  extern virtual task reconfigure_via_task(lvc_configuration cfg);
  extern virtual task wait_for_reset();
  extern task monitor_start();    //monitor start generation
  extern task monitor_stop(lvc_i2c_transaction trans);      //monitor end generation
  extern task ack_counter(logic ack_nack_val);  //count ack/nak number,
  extern task collect_transfer(lvc_i2c_transaction trans);
  extern task data_ana(lvc_i2c_transaction trans);  //analysis collected data from sda line.
  extern task monitor_byte(); // monitor byte unit
  extern task monitor_ack_nack(); // monitor ACK/NACK
  extern task monitor_trans_data(); // monitor byte and ack
  extern function void clear_mon_data();
  extern function void update_trans_data(lvc_i2c_transaction trans); // update trans data from mon_data
endclass

//check all protocol and collect write/read data to transaction
task lvc_i2c_monitor_common::data_ana(lvc_i2c_transaction trans);  
  lvc_i2c_master_transaction mtrans;
  bit addr_first_7bit = 0;
  forever begin
    wait(trans_start_flag | trans_restart_flag);
    trans_restart_flag=0;
    monitor_byte();
    monitor_ack_nack();
    casex(mon_data[mon_data_index])    //check first byte
      8'b0000_001x,8'b0000_010x,8'b0000_011x: begin
        `uvm_error("master monitor common","master monitor receive reserved address")
      end
      8'b0000_0000:  //general call address
      begin
        trans.cmd = I2C_GEN_CALL;
        //collect second byte
        mon_data_index++;
        monitor_byte();
        monitor_ack_nack();
        monitor_trans_data();
        if(trans_restart_flag && mon_data_index!=0) begin
          update_trans_data(trans);
        end
      end
      8'b0000_0001:   //start byte
      begin
        if($cast(mtrans, trans))
          mtrans.send_start_byte = 1'b1;
        trans_start_flag = 0;
        clear_mon_data();
      end
      8'b0000_1xxx:  //hs-mode master code
      begin
        trans_start_flag = 0;
        clear_mon_data();
      end
      8'b1111_1xxx:   //device ID, need check nak and loop.
      begin
        trans.cmd = I2C_DEVICE_ID;
        //devide ID first byte, write slave address followed
        if(mon_data[mon_data_index][0]==0)  begin  
          clear_mon_data();
        end
        //device ID byte followed re-start, read 3 bytes ID
        else if(mon_data[mon_data_index][0]==1)  begin  
          monitor_trans_data();
        end
      end
      8'b1111_0xxx:   //10-bit slave addressing
      begin
        addr_first_7bit = 0;
        if(mon_data[mon_data_index][0]==0)  begin  //10bit address first 7-bits, write
          addr_first_7bit = 1;
          trans.addr_10bit = 1;
          trans.addr[9:8] = mon_data[mon_data_index][2:1];
          mon_data_index++;
          monitor_byte();
          trans.addr[7:0] = mon_data[mon_data_index][7:0];
          monitor_ack_nack();
        end
        if(trans.cmd == I2C_DEVICE_ID) begin
          trans_start_flag = 0;
          clear_mon_data();
        end
        else begin
          trans.cmd = addr_first_7bit ? I2C_WRITE : I2C_READ;
          monitor_trans_data();
          if(trans_restart_flag && mon_data_index != 0) begin
            update_trans_data(trans);
          end
        end
      end
      //normal read and write, should seperate read and write, the last 
      //ack will be a nak generated by master when read.
      default:  
      begin
        if(trans.cmd == I2C_DEVICE_ID) begin
          trans.addr[6:0] = mon_data[mon_data_index][7:1];
          trans_start_flag = 0;
          mon_data = {};
        end
        else begin
          trans.cmd = mon_data[mon_data_index][0] === 0 ? I2C_WRITE : I2C_READ;
          trans.addr[6:0] = mon_data[mon_data_index][7:1];
          monitor_trans_data();
          //10bit address write data with sr end, can sent trans to port
          if(trans_restart_flag && mon_data_index != 0) begin
            update_trans_data(trans);
          end
        end
      end
    endcase
  end
endtask : data_ana

task lvc_i2c_monitor_common::ack_counter(logic ack_nack_val);
  if(ack_nack_val === 0)  //ack
    ack_count++;
  else if(ack_nack_val === 1) //nak
    nack_count++;
  else
    `uvm_error(get_type_name(), $sformatf("ACK_NACK val %b should be 0 or 1", ack_nack_val))
endtask : ack_counter

task lvc_i2c_monitor_common::collect_transfer(lvc_i2c_transaction trans);
  fork
    monitor_start();
    monitor_stop(trans);
    data_ana(trans);
  join_none
endtask : collect_transfer

task lvc_i2c_monitor_common::monitor_start();
  forever begin
    @(negedge i2c_if.SDA);
    begin
      if(i2c_if.SCL == 1 & trans_start_flag == 0) begin
        trans_start_flag = 1;
        trans_stop_flag = 0;
      end
      else if(i2c_if.SCL == 1 & trans_start_flag == 1) begin
        trans_restart_flag = 1;
      end
    end
  end
endtask : monitor_start

task lvc_i2c_monitor_common::monitor_stop(lvc_i2c_transaction trans);
  forever begin
    @(posedge i2c_if.SDA);
    begin
      if(i2c_if.SCL == 1 & trans_start_flag == 1) begin
        update_trans_data(trans);
        trans_stop_flag = 1;
      end
    end
  end
endtask : monitor_stop

task lvc_i2c_monitor_common::monitor_byte(); // monitor byte unit
  for(int i=7;i>=0;i--) begin
    @(posedge i2c_if.SCL);
    mon_data[mon_data_index][i] = i2c_if.SDA;
  end
endtask: monitor_byte

task lvc_i2c_monitor_common::monitor_ack_nack(); 
  logic ack_nack_val;
  @(posedge i2c_if.SCL);
  ack_nack_val = i2c_if.SDA;
  ack_counter(ack_nack_val);
endtask: monitor_ack_nack

task lvc_i2c_monitor_common::monitor_trans_data(); // monitor byte and ack
  logic[8:0] mon_byte; // [8:1] BYTE, [0] ACK/NACK
  logic ack_nack_val;
  int mon_bit_index = 8;
  clear_mon_data();
  while((!trans_stop_flag) & (!trans_restart_flag)) begin
    @(posedge i2c_if.SCL);
    mon_byte[mon_bit_index] = i2c_if.SDA;
    @(negedge i2c_if.SCL);
    if(mon_bit_index==0) begin
      mon_data[mon_data_index] = mon_byte[8:1];
      ack_nack_val = mon_byte[0];
      ack_counter(ack_nack_val);
      mon_bit_index=8;
      mon_data_index++;
    end
    else
      mon_bit_index--;
  end
endtask

function void lvc_i2c_monitor_common::clear_mon_data();
  mon_data_index = 0;
  mon_data = {};
endfunction

function void lvc_i2c_monitor_common::update_trans_data(lvc_i2c_transaction trans); 
  trans.data=mon_data;  
  clear_mon_data();
endfunction

function void lvc_i2c_monitor_common::assign_vif(lvc_i2c_vif i2c_if);
  this.i2c_if = i2c_if;
endfunction

task lvc_i2c_monitor_common::source_event(event sv_e, uvm_event uvm_e);
  forever begin
    @(sv_e);
    uvm_e.trigger();
  end
endtask

task lvc_i2c_monitor_common::reconfigure_via_task(lvc_configuration cfg);
  lvc_i2c_agent_configuration agent_cfg;
  if($cast(agent_cfg,cfg)) begin
    this.cfg.copy(agent_cfg);
  end
  else begin
    `uvm_fatal("CASTFAIL", "I2C configuration handle type inconsistence")
  end
endtask

task lvc_i2c_monitor_common::wait_for_reset();
  // wait for reset release
  @(negedge i2c_if.RST);
endtask

`endif // LVC_I2C_MONITOR_COMMON_SV 
