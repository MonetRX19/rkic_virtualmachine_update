//=======================================================================
// COPYRIGHT (C) 2018-2020 RockerIC, Ltd.
// This software and the associated documentation are confidential and
// proprietary to RockerIC, Ltd. Your use or disclosure of this software
// is subject to the terms and conditions of a consulting agreement
// between you, or your company, and RockerIC, Ltd. In the event of
// publications, the following notice is applicable:
//
// ALL RIGHTS RESERVED
//
// The entire notice above must be reproduced on all authorized copies.
//
// VisitUs  : www.rockeric.com
// Support  : support@rockeric.com
// WeChat   : eva_bill
//-----------------------------------------------------------------------
`ifndef LVC_I2C_DRIVER_COMMON_SV
`define LVC_I2C_DRIVER_COMMON_SV

class lvc_i2c_driver_common extends uvm_object;

  lvc_i2c_vif i2c_if;
  lvc_i2c_agent_configuration cfg;

  `uvm_object_utils_begin(lvc_i2c_driver_common)
  `uvm_object_utils_end
  int unsigned   scl_high_time=0;  //clk high level time
  int unsigned   scl_low_time=0;   //clk low level time
  int unsigned   setup_start_time=0;     //repeat start setup time
  int unsigned   setup_stop_time=0;        //stop setup time
  int unsigned   hold_start_time=0;        //start or repeat start hold time
  int unsigned   hold_data_time=0;        //data hold time
  int unsigned   setup_data_time=0;        //data setup time
  int unsigned   bus_free_time=0;     //bus free time between a stop and start
  int unsigned   data_offset_time=50;   //offset used to sample data for clock strech condition
  bit nack_received_flag = 0;     // flag about nack generated by slave

  extern function new(string name = "lvc_i2c_driver_common");

  extern virtual function void assign_vif(lvc_i2c_vif i2c_if);

  /** source specific event with control variable */
  extern virtual task source_event(event sv_e, uvm_event uvm_e);

  extern virtual task reconfigure_via_task(lvc_configuration cfg);

  //extern virtual task send_xact(lvc_i2c_transaction trans, string type_name);

  //extern virtual task collect_response_from_vif(lvc_i2c_transaction trans);
  extern task wait_data_hold_time(int hold_data_time = this.hold_data_time);
  extern task sda_wait_time_set(int t, logic val);
  extern task scl_wait_time_set(int t, logic val);
  extern task check_slave_ack();
  extern task wait_time(int t);
  extern task extract_time_parameters();
  extern virtual task wait_for_reset();
endclass

function lvc_i2c_driver_common::new(string name = "lvc_i2c_driver_common");
  super.new(name);
endfunction

function void lvc_i2c_driver_common::assign_vif(lvc_i2c_vif i2c_if);
  this.i2c_if = i2c_if;
endfunction

task lvc_i2c_driver_common::source_event(event sv_e, uvm_event uvm_e);
  forever begin
    @(sv_e);
    uvm_e.trigger();
  end
endtask

task lvc_i2c_driver_common::reconfigure_via_task(lvc_configuration cfg);
  lvc_i2c_agent_configuration agent_cfg;

  if($cast(agent_cfg,cfg)) begin
    this.cfg.copy(agent_cfg);
  end
  else begin
    `uvm_fatal("CASTFAIL", "I2C configuration handle type inconsistence")
  end
endtask

task  lvc_i2c_driver_common::extract_time_parameters();
  case (cfg.bus_speed)
    STANDARD_MODE: begin
      scl_high_time    = cfg.scl_high_time_ss;
      scl_low_time     = cfg.scl_low_time_ss;
      setup_start_time = cfg.min_su_sta_time_ss;
      setup_stop_time  = cfg.min_su_sto_time_ss;
      hold_start_time  = cfg.min_hd_sta_time_ss;
      hold_data_time   = cfg.min_hd_dat_time_ss;
      setup_data_time  = cfg.min_su_dat_time_ss;
      bus_free_time    = cfg.tbuf_time_ss;
    end
    FAST_MODE: begin
      scl_high_time    = cfg.scl_high_time_fs;
      scl_low_time     = cfg.scl_low_time_fs;
      setup_start_time = cfg.min_su_sta_time_fs;
      setup_stop_time  = cfg.min_su_sto_time_fs;
      hold_start_time  = cfg.min_hd_sta_time_fs;
      hold_data_time   = cfg.min_hd_dat_time_fs;
      setup_data_time  = cfg.min_su_dat_time_fs;
      bus_free_time    = cfg.tbuf_time_fs;
    end
    HIGHSPEED_MODE: begin
      scl_high_time    = cfg.scl_high_time_hs;
      scl_low_time     = cfg.scl_low_time_hs;
      setup_start_time = cfg.min_su_sta_time_hs;
      setup_stop_time  = cfg.min_su_sto_time_hs;
      hold_start_time  = cfg.min_hd_sta_time_hs;
      hold_data_time   = cfg.min_hd_dat_time_hs;
      setup_data_time  = cfg.min_su_dat_time_hs;
      bus_free_time    = cfg.tbuf_time_hs;
    end
    FAST_MODE_PLUS: begin
      scl_high_time    = cfg.scl_high_time_fm_plus;
      scl_low_time     = cfg.scl_low_time_fm_plus;
      setup_start_time = cfg.min_su_sta_time_fm_plus;
      setup_stop_time  = cfg.min_su_sto_time_fm_plus;
      hold_start_time  = cfg.min_hd_sta_time_fm_plus;
      hold_data_time   = cfg.min_hd_dat_time_fm_plus;
      setup_data_time  = cfg.min_su_dat_time_fm_plus;
      bus_free_time    = cfg.tbuf_time_fm_plus;
    end
    default: begin
      scl_high_time    = cfg.scl_high_time_ss;
      scl_low_time     = cfg.scl_low_time_ss;
      setup_start_time = cfg.min_su_sta_time_ss;
      setup_stop_time  = cfg.min_su_sto_time_ss;
      hold_start_time  = cfg.min_hd_sta_time_ss;
      hold_data_time   = cfg.min_hd_dat_time_ss;
      setup_data_time  = cfg.min_su_dat_time_ss;
      bus_free_time    = cfg.tbuf_time_ss;
    end
  endcase
endtask : extract_time_parameters

task  lvc_i2c_driver_common::wait_data_hold_time(int hold_data_time = this.hold_data_time);
  repeat(hold_data_time) @(posedge i2c_if.CLK);
endtask : wait_data_hold_time

task lvc_i2c_driver_common::wait_time(int t);
  repeat(t) @(posedge i2c_if.CLK);
endtask : wait_time

task lvc_i2c_driver_common::sda_wait_time_set(int t, logic val);
  repeat(t) @(posedge i2c_if.CLK);
  // NOTE:: @Lusang 2020-09-04
  // Use blocking assignment to take effect in case slave drive SDA as
  // 'z' at the same time slot
  i2c_if.sda_master <= val;
endtask : sda_wait_time_set

task lvc_i2c_driver_common::scl_wait_time_set(int t, logic val);
  repeat(t) @(posedge i2c_if.CLK);
  i2c_if.scl_master = val;
  if(val === 1) wait(i2c_if.SCL === val);
endtask : scl_wait_time_set 

task lvc_i2c_driver_common::check_slave_ack();
  if(i2c_if.SDA !=0)
    nack_received_flag = 1;
  else
    nack_received_flag = 0;
endtask: check_slave_ack

task lvc_i2c_driver_common::wait_for_reset();
  // wait for reset release
  @(negedge i2c_if.RST);
endtask

`endif // LVC_I2C_DRIVER_COMMON_SV

